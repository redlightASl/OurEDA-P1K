`timescale 1ns / 1ps 
// `include "linear.v"

module linear_tb();
parameter BITWIDTH = 8;
parameter IS_BITWIDTH_DOUBLE_SCALE = 1;
parameter IN_FEATURES = 14 * 14;
parameter OUT_FEATURES = 10;
parameter USING_BIAS = 0;

reg clk = 0;
reg rst_n = 0;
reg start_sig = 0;

reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_0 = 1568'b11111100_11111000_11010111_11010101_11110011_11110010_11110011_11111001_00000100_00000110_11101000_11010010_11111101_00010010_11101000_11011000_11100000_11110011_11011010_00001001_00001001_00001111_11111101_00010001_00010100_00001100_11110011_00011100_11100110_11101010_11101010_11110100_11110111_11110011_00000101_00000111_11110110_11011110_11011001_11011001_11001100_00100000_11101101_11111000_11110000_11111110_11111100_00001101_00010010_11110110_11011110_11011011_11100101_11000100_11001000_11111001_00000101_00000110_11110100_11111110_11111010_00001110_11011110_11100110_11101100_11101011_11111011_11111011_11100001_11010110_00000010_11111101_11111101_11111100_00000101_11111110_11011111_11010100_11101111_11101100_11111101_00010011_00011001_11111100_00010011_00010100_00011001_00010101_00010011_00001001_11100010_11100110_11111110_00000111_00000110_00010111_00011010_11110001_11110111_00011000_00101000_00101000_00110010_00010110_11011011_11111100_00011110_00001111_00010011_00011001_00101110_00001111_11100100_00000101_00011011_00011100_00110100_00011111_11111010_00000010_00001000_00010001_00001010_00100110_00101011_00101001_11011100_00010101_00011011_00001011_00010011_00010000_11101111_11110110_00001001_00000010_11111110_00000010_00010000_00011100_11100100_00000101_00101110_00010010_00011000_11110110_11110001_00001011_00000100_00000100_11101111_00000001_00000100_00001000_11111101_00011111_11110001_11100001_11001010_10010000_10000000_11010111_00000011_11100011_11101100_11110111_11100111_11111100_11110100_00100000_00100011_11010010_11010000_11000001_11010011_11101011_11001101_11000110_10111000_11001111_11001101_11010111_11101100_11101110_11111101_11110011_11010010_11101011_00000011_00010010_11111000_11111010_11101001_11100001_11011110_11011110;
reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_1 = 1568'b00101001_00110010_10110001_11000111_11111101_11110111_11111100_11011010_11111111_00011010_10111000_10101010_00010011_01001000_11101000_11011110_00100110_00110010_00111001_00101100_00000110_11111110_00000001_00101011_00101010_00011110_11001001_01001100_11011011_11010110_11011001_00101111_01000001_00010110_00101010_00001100_00110110_00110010_00011100_00001000_10111011_00101111_10111111_10111000_10110100_10101011_11011011_11111101_00110111_01000101_00010111_00100111_00011011_00101010_00011101_01010110_11101011_11100001_11000010_10100001_11001010_11111100_00011001_00100101_00011011_00011011_00010101_00011110_00011001_00011011_11101100_00000001_11111101_11010010_11101101_11111011_00001010_00001000_00010111_11101011_11100110_00110001_11101000_11100001_11010010_11101110_11111001_00001111_11100110_00010110_00010011_00001101_00011110_11110000_11011011_11111010_10111110_00001000_10101110_11001000_11001111_11010110_11111011_00010110_00101011_00101000_00101011_00000010_00010100_11010110_11001100_00100111_11010101_11011100_11100111_11011010_00000010_00011101_00110110_00111100_11110110_11101001_11010111_10110011_10000011_11111011_00011000_00100000_00000011_00001011_11101111_00010111_00110111_00110110_11111110_10100100_10100011_11001000_10010111_00001000_00001101_00011010_11111110_11110101_00011001_00110001_00100011_11111000_11001000_10001111_10101000_11010111_11010001_00011000_00000000_00000011_11000001_00010001_11111111_00001100_00000011_11001000_11000101_11010000_00010101_00010101_00001101_00100111_11101110_00010011_00110001_01101010_01111111_00111000_00011010_11111111_11111001_00011101_01000101_00101011_00011101_00100010_10111110_11101000_11100000_00001111_00010000_11111011_10110100_11001011_10111100_11000011_11001101_11010011_11011100_11001100;
reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_2 = 1568'b11111010_11111100_01110110_01111111_01010100_00111110_00111011_00110100_00011000_11100100_11010001_11001111_11101010_11010010_00000101_00011001_00001010_00010011_00001010_11110110_00000110_00010111_11101111_00001100_11110100_11111000_11011101_11100001_00001100_11111001_11101010_11110110_11100000_11100001_11100100_11010111_10111010_10110011_11010011_11110101_00000110_11111110_00010010_00000110_11111100_11111101_00000000_11111011_11101101_11100010_11110010_11100001_11001100_11110010_10110001_00001010_00001000_00000100_00000100_11110111_11010100_11001000_11110011_00010000_00000001_00001111_00010111_00100000_00000010_11010110_11111101_11000111_10101101_10110000_10110101_11011100_00000011_00010001_00100100_00010111_00011000_00100011_00010110_11010110_00011000_11101010_11100000_10101110_11001101_11011010_11111011_00010011_00110000_00110101_00101001_00101001_00100111_00010001_01010000_00001101_11110111_11110000_11101010_11111010_11110100_00000010_00000111_00101110_00011100_00011101_11110110_11111100_01001100_00001000_00010100_00100111_00111001_00010100_11101111_11001001_11011111_11010100_11011110_11000110_11111000_00010010_00001011_00010110_00101011_01000001_00010111_00010010_11100101_11100101_11101001_11001110_11001011_11010000_11000111_00000000_11010110_11100011_00010010_00101100_11111101_00000000_11011101_11101100_11010110_11010001_10110110_11010011_11010011_00001111_11110100_11001010_11100010_11000101_10010110_10010101_10101010_10110110_11000000_11001011_11001100_11101001_11001111_00001001_00010110_00010010_00011100_11100101_11101010_11001011_10011001_10100011_10110011_11100001_11111001_00000011_11111101_00000100_00110010_00110100_01001011_01000011_01000011_00101111_00011100_00001101_11111110_11111000_00000101_00011000_00100010_00101100;
reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_3 = 1568'b00001111_11011011_00001001_11110001_00010010_00010110_00001011_11011100_11011100_11000001_10001010_10000000_11111000_11001110_00101111_11111100_11100111_11100001_00011110_11110111_00001100_00000111_00001101_11101110_11011010_10000011_11010000_11111010_00101111_00001100_11101011_11101101_11100000_11111111_11110111_00000111_11101100_11101100_11100001_10110011_10011010_00011100_00010011_11110011_11010100_11010000_11010111_10111101_10011111_11010001_11100000_11011101_11111001_11110011_00000000_00001111_00001001_11100010_11000111_10111011_10110101_11000110_11111000_00010111_00010001_11111011_11111101_11110110_00010110_00100111_00001000_11001011_10110001_11000100_10110101_11011101_11111100_00001001_00011000_00010001_00010111_00110111_11110101_00001111_00011110_11011110_10111011_11110001_11111000_00001000_00010010_00001000_11100000_00001100_11111111_11111010_00000100_11110111_00100001_11011001_10111100_11100010_11111011_00100010_11101010_11001010_11001001_11001001_11001110_10100100_10101111_11000100_00110100_11111000_11010101_11001011_10111010_11101101_11010010_11010110_11100001_11110101_00001011_11110000_11010100_10100110_00111001_11110110_11011011_11011110_10110001_11011010_11111010_11111100_00010011_00011001_00101101_00010011_00100001_11110001_01000000_00001101_11100010_10111111_10111111_11010010_11010010_11110000_00000100_00010111_00100101_00011011_00101010_00101010_00001010_00101000_00100100_00000111_00000101_11100101_11101011_00001110_00110001_01000100_00100010_00011011_00111000_00101100_11101011_10101001_10010111_10100011_10100110_10110100_11010010_00010011_00100111_00000111_11111011_00001000_00010000_11111100_00011100_00000101_11001011_10001100_10011100_11100000_00000111_00111010_00101011_00110010_01010011_01000100_00111001_01000011;
reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_4 = 1568'b11110111_00010000_10010101_10101101_10101010_11000001_10110011_10110100_10011000_11010011_00100001_00100010_00001011_00101111_00011101_00100110_11111001_11110011_00001100_11011010_11000010_10011010_11001100_11110110_00011000_01000011_00000101_11011101_00011100_00011000_00011111_00011010_00010110_00101001_00000101_00001011_00001111_00010010_00101111_00010011_11111011_11101001_11110001_00011001_00000110_00010010_00011111_00100110_00101100_00111101_01000001_01001100_00010111_11111111_00011100_00001010_11001101_11110001_00000110_00010110_00110100_00110100_00001001_01000001_00110011_00010101_00001101_11110111_00101011_00000001_11100001_00011010_00011100_00010010_00110110_00101010_00101000_00110010_00010001_00011010_00010000_11101010_11111100_00001000_11101100_00000101_00000001_11101111_00000100_11110101_11011001_00000100_00011101_00100101_00010011_11010101_00010010_11100011_11001111_11011010_11110000_11101001_11101111_11001000_10111110_11110100_00000100_00001100_11100101_11111100_11111100_11111010_10101101_11000000_11110110_11110100_11100010_10111101_10111100_11101101_11101011_11101111_11010001_00000011_11000110_11110100_10101000_10000000_10111010_10111110_11011101_11001011_11011111_11011100_11100101_11011011_11110010_11101111_11011010_00000110_11001010_10110000_11100001_00001101_00001000_11101011_11111111_00000111_00000000_11010000_11011100_11010110_11100111_11110111_11101011_00000100_11110111_11111000_00100101_00011110_00110100_00001111_00001001_11110010_11111010_11110011_11110011_11100111_11101010_11111101_00011001_01100011_00111000_00010010_00001111_00010001_00100111_00011000_00101000_00101100_00011100_00000000_11001011_11100111_11111110_00011000_00110100_00010001_11110110_11101100_11001110_11010000_11011101_11100101_11010100_11001011;
reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_5 = 1568'b00000000_11011011_11011110_11001011_11000111_11001101_11100101_11101111_00000100_11101100_11100111_11110100_00010011_00000000_11111011_11111101_00000000_11111010_00000001_11110100_11111011_00001111_00010001_11111001_00001101_00000110_11111001_11011001_00000111_00100110_00010101_00010011_00001001_00000001_00000001_00001010_00010110_00011110_00100101_00100101_00100000_11100011_00000110_00010110_00001111_00001000_00000011_00010001_00010111_00001100_00000111_11110110_11111111_00011010_00001010_00001011_00000100_00000111_00000101_11111100_11111011_00000101_00001011_11001011_11010011_11011110_11011110_11111010_11111000_00010000_00001011_11110101_00000110_00000100_00001111_00000111_11101111_11010011_11000100_11000101_10110100_11001001_11100000_00000100_00010010_11111010_00000011_00000001_00000110_00000010_11110000_11010010_11001010_11000101_10111111_10100111_10100100_11111000_00100000_00001001_11101010_11110001_00000010_00000110_11101001_11100000_11101001_11111010_11100111_11011111_10110111_11110001_00010111_11111001_11100101_11100010_11101011_11110100_11110110_00000011_00000111_11111110_11111001_11101101_00001110_00000011_11111110_11101111_11011100_11100011_11110011_11101110_11111110_00001000_00001101_11111010_00000100_00001000_00001111_00000001_11111000_00000111_11110010_11101100_11101100_11101111_00000111_00001010_11111011_00001101_00010001_00011110_00100101_00000000_11110001_11010011_11110010_11110110_11110111_11111100_00000010_00001011_00010100_00011101_00011000_00100010_00110000_00010101_00010001_11000111_10000000_10101111_11010100_11111100_00000111_11110010_11111111_00000101_00000010_00000111_00000111_00001011_00010111_00011000_11110000_11001110_10111011_11100100_11110010_00000100_00011000_00100011_00010110_00010010_00001111_00010110;
reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_6 = 1568'b11101011_00110100_00111110_00110010_00101001_00100000_00101000_01000100_01111111_01110000_01101011_01011111_11100000_10110101_11101110_00011100_00011000_00001111_11111100_00000110_00001110_00110010_01010001_01000010_00101011_00011011_00101011_00010000_11110101_00010101_00011100_11111100_00001110_11111011_00011100_00001111_00000111_00001010_00001001_00011101_00001100_00101100_11110010_00000011_00100000_00011100_00100100_00100100_00011010_00101111_00001011_00010101_00000100_00010000_00010111_11111100_11110111_00010100_00110111_00101110_00110111_00101011_00001110_00000111_11100101_11010100_11111001_11110111_00010101_00001101_11110111_00101110_00111001_00111001_00110100_00101110_00010011_11110010_10101111_10110001_11000000_11001101_11001110_11010111_11101011_00100111_00101100_00110010_00110110_00011110_00001010_11101011_10101101_10001111_10011011_11011100_11110000_11001001_10111101_00001001_00100000_00011100_00101000_00001110_11111010_11101010_11000111_11010011_11011011_11110011_00001010_00001011_10100101_11110100_00001001_00011101_00110100_00110000_11111001_11101000_11011000_11111101_11110010_00001100_00001010_00000011_10100110_10101000_00011111_00010110_00001111_00001111_00000100_11011001_11101111_11110000_00010001_11110011_11101011_11110110_11011110_11100110_11010010_11100000_00000010_11111000_11010101_11010000_11110001_00001101_00010111_11110011_11011011_11011100_00001100_00100100_11101010_11011100_11010100_10101111_10110100_11010010_11011010_00000000_11110001_11001010_11010111_10110110_11101111_00100110_00100001_10011111_10100101_11011101_11000110_11111011_11110010_11000101_10110110_10110011_10100011_10110000_11101011_11101000_11101101_11111100_11100001_11001111_11110110_11110011_00000111_11111011_11100111_11100100_11010111_11001101;
reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_7 = 1568'b00000001_11110110_11010010_11011011_11001111_11011100_11010111_10110110_10000001_11101000_11011110_11111110_11111011_00001010_00001000_00000100_00001101_11111100_11101010_11011101_11001101_11010110_11001010_11011101_11100110_11011111_11110110_00010110_00010001_00000100_00000000_00000100_11111101_11010110_11100001_11110000_11110000_00000010_11100100_10111010_11011011_00001000_00000111_11111100_11110000_11101010_11100000_11100100_11100110_11111101_00001111_00000110_00010111_11100110_11100101_00000111_11101110_11101111_11101010_11100110_11100101_11001101_11011010_11110100_00001110_11111110_00000100_11110110_11010110_00000101_11111011_11110000_11011100_11111001_11110011_11000110_11001011_11100001_11011110_11111101_00001000_11110010_00000111_11100111_11110100_11110100_11110101_11100100_11101101_00000000_11110111_00001010_00000001_11111001_00000011_11111000_00001101_11100011_11101011_11101110_11110111_11111011_11110011_00000001_00100001_00101010_00011010_00010101_11111110_00000110_00000100_11100001_11011001_11110100_11111100_11111000_11111000_00001101_00000000_00000110_00010101_00100000_00000010_00000101_00001001_00100011_11100111_11011001_11100001_11101101_00010011_00000000_11101101_11111001_11111110_00000000_00000100_00100000_00010111_00101101_00010000_11111011_11110000_00010000_00010100_00010010_00010101_00001010_11110110_11110010_11111100_11110001_11101011_00010000_00000011_00000010_00001001_00001011_00100111_00011110_00010011_00001011_00000110_11110010_11110100_11101111_11010110_11110000_11111100_00010110_00101000_00111100_00100101_00011000_00001101_00010010_00011000_00011100_00001010_11110011_11110011_11101010_11101101_11110110_00010111_00110000_00110100_00010111_00000111_00001000_00010101_00011001_00000010_00000100_11101110_11101110;
reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_8 = 1568'b11111101_11111101_11011111_11101111_11111011_11111110_00010010_00011111_11000110_11000110_11010010_00001111_11110100_11101011_11110111_00000011_00101100_00001110_00011000_00010011_00001011_00001010_11100110_11010001_11101111_11011110_11101000_10100100_11110000_00011011_00011111_00011110_00001000_00011111_00001111_11111010_00011011_11110010_11110101_00110100_01000101_10001110_11111110_00101010_00101001_00101101_00011001_11111010_11000011_10010100_11101011_11101110_00000110_11101010_01010110_10000000_00100001_00000000_00011001_00101110_00000101_00010011_11111010_11001010_00000111_11110011_11010010_00001110_01000000_10110100_11101011_00000111_00010101_00010110_00000101_11100110_00000001_11010100_11110010_00010100_00001001_00011001_01010111_00111110_10110111_11001100_11011101_11011001_11011001_11010010_11101111_11100000_11110010_11101001_00000111_11111101_01000101_01100001_11001011_11110001_11010100_11100000_11011111_11001110_11110111_11101011_00001100_10101100_10100001_11001100_11111100_00011000_11111111_00011111_00101000_00100001_00001001_00010101_00000111_10111010_10010000_10010000_10100110_10110100_11011001_10111000_00001000_01001100_01001100_00111001_01000001_01101011_00011011_11010000_11011101_11100001_11110011_11100001_11110101_11001011_11110110_00010011_00011100_00100011_00100111_00100111_00000101_00001001_00011011_00011000_00010100_00000111_00001000_11010100_11111100_10011100_11010001_00001110_00000101_11010011_10101010_00001001_00100100_00001101_00010111_00001100_00101001_11101101_00110110_00100011_01010101_11000100_10000110_10000101_10001001_11011011_11101110_11100111_11011011_11111011_00001110_11110110_00010111_00011001_00010111_00100001_11000001_10101110_11100001_00000110_00000101_11110000_11110001_00011111_00011011_00100111;
reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_9 = 1568'b11110010_11011011_10101011_11100011_11111010_11011010_11011010_10111001_11101111_10110011_10000000_11101010_11110110_00010000_11011000_11010110_11010011_11011010_11110001_00010001_11110110_00011110_00101110_11111100_10111010_11100001_00000000_00101110_11010111_11100011_11100110_11011110_11101111_00000101_11111100_11111010_00000101_00001100_11001111_10100001_11010011_00000100_00000111_11111000_00001110_00011011_00010000_11100110_11010010_11000101_11001001_11001010_11000010_10110011_10110101_00001010_00100011_00100011_00101000_00100111_00011111_00001011_11101100_11011001_11010000_11100100_11100010_11010101_11011111_00010010_00010001_00100000_00010000_00010001_11111101_00000011_11101101_00010100_00001011_00000101_00010000_11110010_11011001_00010001_11110110_00001011_00001100_00010000_11111010_11011001_00001001_11111111_00000101_11111100_00010001_11111100_11000001_00001111_11011001_00000110_00010000_00000110_11011110_10111011_11101100_00000100_00000100_11111100_00010100_00010000_11111010_00100010_11100110_00000110_11110111_11110110_10110100_10011011_11100000_11111001_00011000_00000111_00000011_11101101_11101100_11100110_11111111_00001010_11111000_11101000_11001000_11010000_00000111_00000010_00010001_00001111_11111011_11101010_11010011_11000001_00010110_00100101_11101111_11101111_11010001_11111100_00001011_00010001_00001111_11111011_11111110_00000000_00001000_11001111_00010101_01000000_00100101_00000101_00001101_00101000_00100110_00100110_11111110_11111001_11110000_11101001_11101000_11101001_00000100_00010011_11111001_11101100_00001111_00100011_00010101_00000001_11110111_11111000_11111010_11111111_00010000_00111110_11111001_00000101_11110011_11111001_00010001_00011101_00010110_11110110_11110110_11111011_11111001_11111000_11100111_11101111;

// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_9 = 1568'b11111100_11111000_11010111_11010101_11110011_11110010_11110011_11111001_00000100_00000110_11101000_11010010_11111101_00010010_11101000_11011000_11100000_11110011_11011010_00001001_00001001_00001111_11111101_00010001_00010100_00001100_11110011_00011100_11100110_11101010_11101010_11110100_11110111_11110011_00000101_00000111_11110110_11011110_11011001_11011001_11001100_00100000_11101101_11111000_11110000_11111110_11111100_00001101_00010010_11110110_11011110_11011011_11100101_11000100_11001000_11111001_00000101_00000110_11110100_11111110_11111010_00001110_11011110_11100110_11101100_11101011_11111011_11111011_11100001_11010110_00000010_11111101_11111101_11111100_00000101_11111110_11011111_11010100_11101111_11101100_11111101_00010011_00011001_11111100_00010011_00010100_00011001_00010101_00010011_00001001_11100010_11100110_11111110_00000111_00000110_00010111_00011010_11110001_11110111_00011000_00101000_00101000_00110010_00010110_11011011_11111100_00011110_00001111_00010011_00011001_00101110_00001111_11100100_00000101_00011011_00011100_00110100_00011111_11111010_00000010_00001000_00010001_00001010_00100110_00101011_00101001_11011100_00010101_00011011_00001011_00010011_00010000_11101111_11110110_00001001_00000010_11111110_00000010_00010000_00011100_11100100_00000101_00101110_00010010_00011000_11110110_11110001_00001011_00000100_00000100_11101111_00000001_00000100_00001000_11111101_00011111_11110001_11100001_11001010_10010000_10000000_11010111_00000011_11100011_11101100_11110111_11100111_11111100_11110100_00100000_00100011_11010010_11010000_11000001_11010011_11101011_11001101_11000110_10111000_11001111_11001101_11010111_11101100_11101110_11111101_11110011_11010010_11101011_00000011_00010010_11111000_11111010_11101001_11100001_11011110_11011110;
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_8 = 1568'b00101001_00110010_10110001_11000111_11111101_11110111_11111100_11011010_11111111_00011010_10111000_10101010_00010011_01001000_11101000_11011110_00100110_00110010_00111001_00101100_00000110_11111110_00000001_00101011_00101010_00011110_11001001_01001100_11011011_11010110_11011001_00101111_01000001_00010110_00101010_00001100_00110110_00110010_00011100_00001000_10111011_00101111_10111111_10111000_10110100_10101011_11011011_11111101_00110111_01000101_00010111_00100111_00011011_00101010_00011101_01010110_11101011_11100001_11000010_10100001_11001010_11111100_00011001_00100101_00011011_00011011_00010101_00011110_00011001_00011011_11101100_00000001_11111101_11010010_11101101_11111011_00001010_00001000_00010111_11101011_11100110_00110001_11101000_11100001_11010010_11101110_11111001_00001111_11100110_00010110_00010011_00001101_00011110_11110000_11011011_11111010_10111110_00001000_10101110_11001000_11001111_11010110_11111011_00010110_00101011_00101000_00101011_00000010_00010100_11010110_11001100_00100111_11010101_11011100_11100111_11011010_00000010_00011101_00110110_00111100_11110110_11101001_11010111_10110011_10000011_11111011_00011000_00100000_00000011_00001011_11101111_00010111_00110111_00110110_11111110_10100100_10100011_11001000_10010111_00001000_00001101_00011010_11111110_11110101_00011001_00110001_00100011_11111000_11001000_10001111_10101000_11010111_11010001_00011000_00000000_00000011_11000001_00010001_11111111_00001100_00000011_11001000_11000101_11010000_00010101_00010101_00001101_00100111_11101110_00010011_00110001_01101010_01111111_00111000_00011010_11111111_11111001_00011101_01000101_00101011_00011101_00100010_10111110_11101000_11100000_00001111_00010000_11111011_10110100_11001011_10111100_11000011_11001101_11010011_11011100_11001100;
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_7 = 1568'b11111010_11111100_01110110_01111111_01010100_00111110_00111011_00110100_00011000_11100100_11010001_11001111_11101010_11010010_00000101_00011001_00001010_00010011_00001010_11110110_00000110_00010111_11101111_00001100_11110100_11111000_11011101_11100001_00001100_11111001_11101010_11110110_11100000_11100001_11100100_11010111_10111010_10110011_11010011_11110101_00000110_11111110_00010010_00000110_11111100_11111101_00000000_11111011_11101101_11100010_11110010_11100001_11001100_11110010_10110001_00001010_00001000_00000100_00000100_11110111_11010100_11001000_11110011_00010000_00000001_00001111_00010111_00100000_00000010_11010110_11111101_11000111_10101101_10110000_10110101_11011100_00000011_00010001_00100100_00010111_00011000_00100011_00010110_11010110_00011000_11101010_11100000_10101110_11001101_11011010_11111011_00010011_00110000_00110101_00101001_00101001_00100111_00010001_01010000_00001101_11110111_11110000_11101010_11111010_11110100_00000010_00000111_00101110_00011100_00011101_11110110_11111100_01001100_00001000_00010100_00100111_00111001_00010100_11101111_11001001_11011111_11010100_11011110_11000110_11111000_00010010_00001011_00010110_00101011_01000001_00010111_00010010_11100101_11100101_11101001_11001110_11001011_11010000_11000111_00000000_11010110_11100011_00010010_00101100_11111101_00000000_11011101_11101100_11010110_11010001_10110110_11010011_11010011_00001111_11110100_11001010_11100010_11000101_10010110_10010101_10101010_10110110_11000000_11001011_11001100_11101001_11001111_00001001_00010110_00010010_00011100_11100101_11101010_11001011_10011001_10100011_10110011_11100001_11111001_00000011_11111101_00000100_00110010_00110100_01001011_01000011_01000011_00101111_00011100_00001101_11111110_11111000_00000101_00011000_00100010_00101100;
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_6 = 1568'b00001111_11011011_00001001_11110001_00010010_00010110_00001011_11011100_11011100_11000001_10001010_10000000_11111000_11001110_00101111_11111100_11100111_11100001_00011110_11110111_00001100_00000111_00001101_11101110_11011010_10000011_11010000_11111010_00101111_00001100_11101011_11101101_11100000_11111111_11110111_00000111_11101100_11101100_11100001_10110011_10011010_00011100_00010011_11110011_11010100_11010000_11010111_10111101_10011111_11010001_11100000_11011101_11111001_11110011_00000000_00001111_00001001_11100010_11000111_10111011_10110101_11000110_11111000_00010111_00010001_11111011_11111101_11110110_00010110_00100111_00001000_11001011_10110001_11000100_10110101_11011101_11111100_00001001_00011000_00010001_00010111_00110111_11110101_00001111_00011110_11011110_10111011_11110001_11111000_00001000_00010010_00001000_11100000_00001100_11111111_11111010_00000100_11110111_00100001_11011001_10111100_11100010_11111011_00100010_11101010_11001010_11001001_11001001_11001110_10100100_10101111_11000100_00110100_11111000_11010101_11001011_10111010_11101101_11010010_11010110_11100001_11110101_00001011_11110000_11010100_10100110_00111001_11110110_11011011_11011110_10110001_11011010_11111010_11111100_00010011_00011001_00101101_00010011_00100001_11110001_01000000_00001101_11100010_10111111_10111111_11010010_11010010_11110000_00000100_00010111_00100101_00011011_00101010_00101010_00001010_00101000_00100100_00000111_00000101_11100101_11101011_00001110_00110001_01000100_00100010_00011011_00111000_00101100_11101011_10101001_10010111_10100011_10100110_10110100_11010010_00010011_00100111_00000111_11111011_00001000_00010000_11111100_00011100_00000101_11001011_10001100_10011100_11100000_00000111_00111010_00101011_00110010_01010011_01000100_00111001_01000011;
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_5 = 1568'b11110111_00010000_10010101_10101101_10101010_11000001_10110011_10110100_10011000_11010011_00100001_00100010_00001011_00101111_00011101_00100110_11111001_11110011_00001100_11011010_11000010_10011010_11001100_11110110_00011000_01000011_00000101_11011101_00011100_00011000_00011111_00011010_00010110_00101001_00000101_00001011_00001111_00010010_00101111_00010011_11111011_11101001_11110001_00011001_00000110_00010010_00011111_00100110_00101100_00111101_01000001_01001100_00010111_11111111_00011100_00001010_11001101_11110001_00000110_00010110_00110100_00110100_00001001_01000001_00110011_00010101_00001101_11110111_00101011_00000001_11100001_00011010_00011100_00010010_00110110_00101010_00101000_00110010_00010001_00011010_00010000_11101010_11111100_00001000_11101100_00000101_00000001_11101111_00000100_11110101_11011001_00000100_00011101_00100101_00010011_11010101_00010010_11100011_11001111_11011010_11110000_11101001_11101111_11001000_10111110_11110100_00000100_00001100_11100101_11111100_11111100_11111010_10101101_11000000_11110110_11110100_11100010_10111101_10111100_11101101_11101011_11101111_11010001_00000011_11000110_11110100_10101000_10000000_10111010_10111110_11011101_11001011_11011111_11011100_11100101_11011011_11110010_11101111_11011010_00000110_11001010_10110000_11100001_00001101_00001000_11101011_11111111_00000111_00000000_11010000_11011100_11010110_11100111_11110111_11101011_00000100_11110111_11111000_00100101_00011110_00110100_00001111_00001001_11110010_11111010_11110011_11110011_11100111_11101010_11111101_00011001_01100011_00111000_00010010_00001111_00010001_00100111_00011000_00101000_00101100_00011100_00000000_11001011_11100111_11111110_00011000_00110100_00010001_11110110_11101100_11001110_11010000_11011101_11100101_11010100_11001011;
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_4 = 1568'b00000000_11011011_11011110_11001011_11000111_11001101_11100101_11101111_00000100_11101100_11100111_11110100_00010011_00000000_11111011_11111101_00000000_11111010_00000001_11110100_11111011_00001111_00010001_11111001_00001101_00000110_11111001_11011001_00000111_00100110_00010101_00010011_00001001_00000001_00000001_00001010_00010110_00011110_00100101_00100101_00100000_11100011_00000110_00010110_00001111_00001000_00000011_00010001_00010111_00001100_00000111_11110110_11111111_00011010_00001010_00001011_00000100_00000111_00000101_11111100_11111011_00000101_00001011_11001011_11010011_11011110_11011110_11111010_11111000_00010000_00001011_11110101_00000110_00000100_00001111_00000111_11101111_11010011_11000100_11000101_10110100_11001001_11100000_00000100_00010010_11111010_00000011_00000001_00000110_00000010_11110000_11010010_11001010_11000101_10111111_10100111_10100100_11111000_00100000_00001001_11101010_11110001_00000010_00000110_11101001_11100000_11101001_11111010_11100111_11011111_10110111_11110001_00010111_11111001_11100101_11100010_11101011_11110100_11110110_00000011_00000111_11111110_11111001_11101101_00001110_00000011_11111110_11101111_11011100_11100011_11110011_11101110_11111110_00001000_00001101_11111010_00000100_00001000_00001111_00000001_11111000_00000111_11110010_11101100_11101100_11101111_00000111_00001010_11111011_00001101_00010001_00011110_00100101_00000000_11110001_11010011_11110010_11110110_11110111_11111100_00000010_00001011_00010100_00011101_00011000_00100010_00110000_00010101_00010001_11000111_10000000_10101111_11010100_11111100_00000111_11110010_11111111_00000101_00000010_00000111_00000111_00001011_00010111_00011000_11110000_11001110_10111011_11100100_11110010_00000100_00011000_00100011_00010110_00010010_00001111_00010110;
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_3 = 1568'b11101011_00110100_00111110_00110010_00101001_00100000_00101000_01000100_01111111_01110000_01101011_01011111_11100000_10110101_11101110_00011100_00011000_00001111_11111100_00000110_00001110_00110010_01010001_01000010_00101011_00011011_00101011_00010000_11110101_00010101_00011100_11111100_00001110_11111011_00011100_00001111_00000111_00001010_00001001_00011101_00001100_00101100_11110010_00000011_00100000_00011100_00100100_00100100_00011010_00101111_00001011_00010101_00000100_00010000_00010111_11111100_11110111_00010100_00110111_00101110_00110111_00101011_00001110_00000111_11100101_11010100_11111001_11110111_00010101_00001101_11110111_00101110_00111001_00111001_00110100_00101110_00010011_11110010_10101111_10110001_11000000_11001101_11001110_11010111_11101011_00100111_00101100_00110010_00110110_00011110_00001010_11101011_10101101_10001111_10011011_11011100_11110000_11001001_10111101_00001001_00100000_00011100_00101000_00001110_11111010_11101010_11000111_11010011_11011011_11110011_00001010_00001011_10100101_11110100_00001001_00011101_00110100_00110000_11111001_11101000_11011000_11111101_11110010_00001100_00001010_00000011_10100110_10101000_00011111_00010110_00001111_00001111_00000100_11011001_11101111_11110000_00010001_11110011_11101011_11110110_11011110_11100110_11010010_11100000_00000010_11111000_11010101_11010000_11110001_00001101_00010111_11110011_11011011_11011100_00001100_00100100_11101010_11011100_11010100_10101111_10110100_11010010_11011010_00000000_11110001_11001010_11010111_10110110_11101111_00100110_00100001_10011111_10100101_11011101_11000110_11111011_11110010_11000101_10110110_10110011_10100011_10110000_11101011_11101000_11101101_11111100_11100001_11001111_11110110_11110011_00000111_11111011_11100111_11100100_11010111_11001101;
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_2 = 1568'b00000001_11110110_11010010_11011011_11001111_11011100_11010111_10110110_10000001_11101000_11011110_11111110_11111011_00001010_00001000_00000100_00001101_11111100_11101010_11011101_11001101_11010110_11001010_11011101_11100110_11011111_11110110_00010110_00010001_00000100_00000000_00000100_11111101_11010110_11100001_11110000_11110000_00000010_11100100_10111010_11011011_00001000_00000111_11111100_11110000_11101010_11100000_11100100_11100110_11111101_00001111_00000110_00010111_11100110_11100101_00000111_11101110_11101111_11101010_11100110_11100101_11001101_11011010_11110100_00001110_11111110_00000100_11110110_11010110_00000101_11111011_11110000_11011100_11111001_11110011_11000110_11001011_11100001_11011110_11111101_00001000_11110010_00000111_11100111_11110100_11110100_11110101_11100100_11101101_00000000_11110111_00001010_00000001_11111001_00000011_11111000_00001101_11100011_11101011_11101110_11110111_11111011_11110011_00000001_00100001_00101010_00011010_00010101_11111110_00000110_00000100_11100001_11011001_11110100_11111100_11111000_11111000_00001101_00000000_00000110_00010101_00100000_00000010_00000101_00001001_00100011_11100111_11011001_11100001_11101101_00010011_00000000_11101101_11111001_11111110_00000000_00000100_00100000_00010111_00101101_00010000_11111011_11110000_00010000_00010100_00010010_00010101_00001010_11110110_11110010_11111100_11110001_11101011_00010000_00000011_00000010_00001001_00001011_00100111_00011110_00010011_00001011_00000110_11110010_11110100_11101111_11010110_11110000_11111100_00010110_00101000_00111100_00100101_00011000_00001101_00010010_00011000_00011100_00001010_11110011_11110011_11101010_11101101_11110110_00010111_00110000_00110100_00010111_00000111_00001000_00010101_00011001_00000010_00000100_11101110_11101110;
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_1 = 1568'b11111101_11111101_11011111_11101111_11111011_11111110_00010010_00011111_11000110_11000110_11010010_00001111_11110100_11101011_11110111_00000011_00101100_00001110_00011000_00010011_00001011_00001010_11100110_11010001_11101111_11011110_11101000_10100100_11110000_00011011_00011111_00011110_00001000_00011111_00001111_11111010_00011011_11110010_11110101_00110100_01000101_10001110_11111110_00101010_00101001_00101101_00011001_11111010_11000011_10010100_11101011_11101110_00000110_11101010_01010110_10000000_00100001_00000000_00011001_00101110_00000101_00010011_11111010_11001010_00000111_11110011_11010010_00001110_01000000_10110100_11101011_00000111_00010101_00010110_00000101_11100110_00000001_11010100_11110010_00010100_00001001_00011001_01010111_00111110_10110111_11001100_11011101_11011001_11011001_11010010_11101111_11100000_11110010_11101001_00000111_11111101_01000101_01100001_11001011_11110001_11010100_11100000_11011111_11001110_11110111_11101011_00001100_10101100_10100001_11001100_11111100_00011000_11111111_00011111_00101000_00100001_00001001_00010101_00000111_10111010_10010000_10010000_10100110_10110100_11011001_10111000_00001000_01001100_01001100_00111001_01000001_01101011_00011011_11010000_11011101_11100001_11110011_11100001_11110101_11001011_11110110_00010011_00011100_00100011_00100111_00100111_00000101_00001001_00011011_00011000_00010100_00000111_00001000_11010100_11111100_10011100_11010001_00001110_00000101_11010011_10101010_00001001_00100100_00001101_00010111_00001100_00101001_11101101_00110110_00100011_01010101_11000100_10000110_10000101_10001001_11011011_11101110_11100111_11011011_11111011_00001110_11110110_00010111_00011001_00010111_00100001_11000001_10101110_11100001_00000110_00000101_11110000_11110001_00011111_00011011_00100111;
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_0 = 1568'b11110010_11011011_10101011_11100011_11111010_11011010_11011010_10111001_11101111_10110011_10000000_11101010_11110110_00010000_11011000_11010110_11010011_11011010_11110001_00010001_11110110_00011110_00101110_11111100_10111010_11100001_00000000_00101110_11010111_11100011_11100110_11011110_11101111_00000101_11111100_11111010_00000101_00001100_11001111_10100001_11010011_00000100_00000111_11111000_00001110_00011011_00010000_11100110_11010010_11000101_11001001_11001010_11000010_10110011_10110101_00001010_00100011_00100011_00101000_00100111_00011111_00001011_11101100_11011001_11010000_11100100_11100010_11010101_11011111_00010010_00010001_00100000_00010000_00010001_11111101_00000011_11101101_00010100_00001011_00000101_00010000_11110010_11011001_00010001_11110110_00001011_00001100_00010000_11111010_11011001_00001001_11111111_00000101_11111100_00010001_11111100_11000001_00001111_11011001_00000110_00010000_00000110_11011110_10111011_11101100_00000100_00000100_11111100_00010100_00010000_11111010_00100010_11100110_00000110_11110111_11110110_10110100_10011011_11100000_11111001_00011000_00000111_00000011_11101101_11101100_11100110_11111111_00001010_11111000_11101000_11001000_11010000_00000111_00000010_00010001_00001111_11111011_11101010_11010011_11000001_00010110_00100101_11101111_11101111_11010001_11111100_00001011_00010001_00001111_11111011_11111110_00000000_00001000_11001111_00010101_01000000_00100101_00000101_00001101_00101000_00100110_00100110_11111110_11111001_11110000_11101001_11101000_11101001_00000100_00010011_11111001_11101100_00001111_00100011_00010101_00000001_11110111_11111000_11111010_11111111_00010000_00111110_11111001_00000101_11110011_11111001_00010001_00011101_00010110_11110110_11110110_11111011_11111001_11111000_11100111_11101111;

// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_0 = {14*14{8'b0000_0001}};
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_1 = {14*14{8'b0000_0001}};
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_2 = {14*14{8'b0000_0001}};
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_3 = {14*14{8'b0000_0001}};
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_4 = {14*14{8'b0000_0001}};
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_5 = {14*14{8'b0000_0001}};
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_6 = {14*14{8'b0000_0001}};
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_7 = {14*14{8'b0000_0001}};
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_8 = {14*14{8'b0000_0001}};
// reg signed [IN_FEATURES * BITWIDTH - 1 : 0] weight_mem_9 = {14*14{8'b0000_0001}};

reg signed [OUT_FEATURES * BITWIDTH * (IS_BITWIDTH_DOUBLE_SCALE + 1) - 1 : 0] bias_mem = {(OUT_FEATURES * BITWIDTH * (IS_BITWIDTH_DOUBLE_SCALE + 1)){1'b0}};
reg signed [BITWIDTH * IN_FEATURES - 1 : 0] in_features = 1568'b0;

// linear Outputs
wire signed [BITWIDTH * (IS_BITWIDTH_DOUBLE_SCALE + 1) * OUT_FEATURES - 1 : 0] out_features;

wire [BITWIDTH - 1: 0] output_data_0;
wire [BITWIDTH - 1: 0] output_data_1;
wire [BITWIDTH - 1: 0] output_data_2;
wire [BITWIDTH - 1: 0] output_data_3;
wire [BITWIDTH - 1: 0] output_data_4;
wire [BITWIDTH - 1: 0] output_data_5;
wire [BITWIDTH - 1: 0] output_data_6;
wire [BITWIDTH - 1: 0] output_data_7;
wire [BITWIDTH - 1: 0] output_data_8;
wire [BITWIDTH - 1: 0] output_data_9;

// assign {output_data_0, output_data_1, output_data_2, output_data_3, output_data_4, output_data_5, output_data_6, output_data_7, output_data_8, output_data_9} = out_features;
assign output_data_9 = out_features[7:0];
assign output_data_8 = out_features[23:16];
assign output_data_7 = out_features[39:32];
assign output_data_6 = out_features[55:48];
assign output_data_5 = out_features[71:64];
assign output_data_4 = out_features[87:80];
assign output_data_3 = out_features[103:96];
assign output_data_2 = out_features[119:112];
assign output_data_1 = out_features[135:128];
assign output_data_0 = out_features[151:144];

wire done_sig;

initial begin
    forever
        #5 clk = ~clk;
end

/*
weight=正常
data=全1
-81,  31, -95, -90, -93, -43,  83,  77, -56,  20
00AF 001F 00A1 00A6 00A3 00D5 0053 004D 00C8 0014
*/

/*
weight=全1
data=全1
-60, -60, -60, -60, -60, -60, -60, -60, -60, -60
C4 C4 C4 C4 C4 C4 C4 C4 C4 C4
*/


integer stage = 0;
always @(posedge clk) begin
    case (stage)
        0: begin
            rst_n = 1'b1;
            start_sig = 1'b0;
            stage = 1;
        end
        1: begin
            in_features = {14 * 14{8'b0000_0101}};
            // in_features = {1568{1'b0}};
            start_sig = 1'b1;
            stage = 2;
        end
        2: begin
            stage = 3;
        end
        3: begin
            stage = 4;
        end
        4: begin
            if (done_sig) begin
                in_features <= {1568{1'b0}};
                weight_mem_0 <= {1568{1'b0}};
                weight_mem_1 <= {1568{1'b0}};
                weight_mem_2 <= {1568{1'b0}};
                weight_mem_3 <= {1568{1'b0}};
                weight_mem_4 <= {1568{1'b0}};
                weight_mem_5 <= {1568{1'b0}};
                weight_mem_6 <= {1568{1'b0}};
                weight_mem_7 <= {1568{1'b0}};
                weight_mem_8 <= {1568{1'b0}};
                weight_mem_9 <= {1568{1'b0}};
                start_sig = 1'b0;
                stage = 5;
                $display("%d", $signed(output_data_0));
                $display("%d", $signed(output_data_1));
                $display("%d", $signed(output_data_2));
                $display("%d", $signed(output_data_3));
                $display("%d", $signed(output_data_4));
                $display("%d", $signed(output_data_5));
                $display("%d", $signed(output_data_6));
                $display("%d", $signed(output_data_7));
                $display("%d", $signed(output_data_8));
                $display("%d", $signed(output_data_9));
                // $display("%b",output_data_0);
                // $display("%d",output_data_1);
                // $display("%d",output_data_2);
                // $display("%d",output_data_3);
                // $display("%d",output_data_4);
                // $display("%d",output_data_5);
                // $display("%d",output_data_6);
                // $display("%d",output_data_7);
                // $display("%d",output_data_8);
                // $display("%d",output_data_9);
            end
            else begin
                stage = 4;
            end
        end
        default: begin

        end
    endcase
end


initial begin
    $dumpfile("linear_tb.vcd");
    $dumpvars();
    #500;
    #500;
    #500;
    #500;
    #500;
    #500;
    #500;
    #500;
    #500;
    #500;
    $finish;
end

linear #(
           .BITWIDTH ( BITWIDTH ),
           .IS_BITWIDTH_DOUBLE_SCALE( IS_BITWIDTH_DOUBLE_SCALE ),
           .IN_FEATURES ( IN_FEATURES ),
           .OUT_FEATURES ( OUT_FEATURES ),
           .USING_BIAS ( USING_BIAS ))
       u_linear(
           //ports
           .clk ( clk ),
           .rst_n ( rst_n ),
           .valid ( start_sig ),
           .ready ( done_sig ),
           .weight_mem_0 ( weight_mem_0 ),
           .weight_mem_1 ( weight_mem_1 ),
           .weight_mem_2 ( weight_mem_2 ),
           .weight_mem_3 ( weight_mem_3 ),
           .weight_mem_4 ( weight_mem_4 ),
           .weight_mem_5 ( weight_mem_5 ),
           .weight_mem_6 ( weight_mem_6 ),
           .weight_mem_7 ( weight_mem_7 ),
           .weight_mem_8 ( weight_mem_8 ),
           .weight_mem_9 ( weight_mem_9 ),
           .bias_mem ( bias_mem ),
           .in_features ( in_features ),
           .out_features ( out_features )
       );

endmodule

